<?xml version="1.0" encoding="UTF-8"?>
<Batch version="1.0"><TaskList><Task type="ResizeTask" enabled="True"><Width units="0">4000</Width><Height units="0">-1</Height><DPI>-1</DPI><Filter>9</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType></Task></TaskList></Batch>
